`include "CLA8.v"

module CLA32(
    input  [31:0] a,
    input  [31:0] b,
    output [31:0] sum,
    output overflow);

// put your design here

endmodule