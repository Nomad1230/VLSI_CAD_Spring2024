module black_cell(p1, p2, g1, g2, G, P);
input  p1, p2, g1, g2;
output G, P;

// put your design here

endmodule