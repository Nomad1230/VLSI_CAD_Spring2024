module FA(
    input  a,
    input  b,
    input  Cin, 
    output Sum,
    output cout);

// put your design here

endmodule