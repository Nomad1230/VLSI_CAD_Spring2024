`include "RCA4.v"

module RCA16(
    input  [15:0] a,
    input  [15:0] b,
    output [15:0] sum,
    output overflow
);

// put your design here

endmodule