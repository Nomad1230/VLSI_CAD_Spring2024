module FA(
    input  a,
    input  b,
    input  cin, 
    output sum,
    output cout
);

	// put your design here

endmodule