`include "black_cell.v"
`include "blue_cell.v"

module PPA8(A, B, Cin, Sum, Cout);
input  [7:0] A, B;
input        Cin;
output [7:0] Sum;
output Cout;

// put your design here


endmodule