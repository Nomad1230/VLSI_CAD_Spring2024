// ================================================ // 
//  Course:      IVCAD 2024 Spring                  //                       
//  Auther:      Zong-Jin CAI (Leo)                 //                         
//  Filename:    Multiplier_PPA.v                   //                               
//  Description: 8*8-bit Multiplier using PPA       //                 
//  Version:     1.0                                // 
//  Date:        2024/02/22                         //     
// ================================================ //    

`include "PPA8.v"

module Multiplier_PPA(
    input   [7:0]   A,
    input   [7:0]   B,
    output  [15:0]  Product
);
    // put your design here
    
endmodule
