module blue_cell(p2, g1, g2, G);
input  p2, g1, g2;
output G;

// put your design here

endmodule