// ================================================ // 
//  Course:      IVCAD 2024 Spring                  //                       
//  Auther:      Zong-Jin CAI (Leo)                 //                         
//  Filename:    PPA.v                              //                               
//  Description: Parallel Prefix Adder              //                 
//  Version:     1.0                                // 
//  Date:        2024/02/22                         //     
//  Reference:   Yong-Sheng Liu (David)             //
// ================================================ //   
`include "black_cell.v"
`include "blue_cell.v"

module PPA8(A, B, Cin, Sum, Cout);
input  [7:0] A, B;
input        Cin;
output [7:0] Sum;
output Cout;

// put your design here

endmodule